`default_nettype none

/* verilator lint_off UNUSED */

module tt_um_urish_simon (
	input  wire [7:0] ui_in,	// Dedicated inputs
	output wire [7:0] uo_out,	// Dedicated outputs
	input  wire [7:0] uio_in,	// IOs: Input path
	output wire [7:0] uio_out,	// IOs: Output path
	output wire [7:0] uio_oe,	// IOs: Enable path (active high: 0=input, 1=output)
	input  wire       ena,
	input  wire       clk,
	input  wire       rst_n
);

  wire [3:0]led;
  wire sound;

  assign uo_out = { 3'b0, sound, led };
  assign uio_oe = 0;
  assign uio_out = 0;

  simon simon1 (
      .clk   (clk),
      .rst   (!rst_n),
      .ticks_per_milli (50),
      .btn   (ui_in[3:0]),
      .led   (led),
      .sound (sound)
  );

endmodule
